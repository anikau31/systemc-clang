module sreg_0(
  input clk,
  input reset
);

endmodule // sreg_0

module sreg_1(
  input clk,
  input reset
);

endmodule // sreg_1

module sreg_2(
  input clk,
  input reset
);

endmodule // sreg_2
