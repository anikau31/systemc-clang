program automatic test_case(); // interface to the design
  initial begin
    $display("Test case");
  end
endprogram


